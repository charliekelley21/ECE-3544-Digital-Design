////////////////////////////////////////////////////////////////////////////////
// Filename:    tb_project3a.v
// Author:      J.S. Thweatt
// Date:        08 October 2015
// Version:     1
// Description: This is the skeleton of a test bench for Project 3A. UPDATE
//              THIS DESCRIPTION WHEN YOU IMPLEMENT YOUR TEST BENCH.

`timescale 1 ns/100 ps

module tb_project3a();
//  Declare regs and wires.



//  Instantiate system.



//  Test the circuit functionality here. You should apply different combinations
//  of the inputs and observer the outputs for correctness.



//  This is not the only module that you could have tested. As long as you can
//  write a test bench, add it to your project, and follow the instructions for
//  invoking ModelSim from Quartus, you can test any module that you create in
//  Quartus.

endmodule
