// DELETE THESE COMMENTS AFTER YOU ADD YOUR MODULE HEADER HERE.
// Insert a module header in the style of the starter code and review module on Verilog fundamentals.
// Your description should include your input assignment.

// DELETE THESE COMMENTS AFTER YOU RENAME YOUR FILE AND ADD IT TO THE PROJECT
// Insert your Virginia Tech PID into part of the module name labeled YOURPID.
// - Your Virginia Tech PID is the part of your e-mail address preceding "@vt.edu".
// Save your file with the complete name of your module, then add the re-named file to the project.
// - Right-click in the Project Window, choose Add to Project > Existing File, then Browse for the file.
// Remove the original file from the Project. You don't have to delete the file from your disk.
// - Right-click the file name in the Project Window, and choose Remove from Project.

module rpsJudge_structural_YOURPID(player1, player2, p1wins, p2wins, tied);
   input  [2:0] player1, player2;
   output       p1wins, p2wins, tied;

   // Your module MUST consist solely of primitive logic gates.
   // Declare additional wires as needed.


endmodule
